
`ifndef MODULE_PARAMETER
    `define ROB_DEPTH 8
    `define DATA_WIDTH 32
`endif
